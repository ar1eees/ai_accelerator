module top_streaming_acc (
    input clk, nrst, 
);
    
endmodule